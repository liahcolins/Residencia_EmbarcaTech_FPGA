module porta_not(
    input logic a,
    output logic y
);

    assign y = ~a;
endmodule